initial begin
    $readmemh("softplus_lut.mem", lut_mem);
end
